//
// Verilog Module cat_recognizer_lib.stimulus_direct
//
// Created:
//          by - amitb.UNKNOWN (DESKTOP-GIFQ7HQ)
//          at - 13:32:43 15/12/2018
//
// using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
//

`resetall
`timescale 1ns/10ps
module stimulus_direct ;


// ### Please start your Verilog code here ### 

endmodule
