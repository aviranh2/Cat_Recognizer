//
// Verilog Module cat_recognizer_lib.checker
//
// Created:
//          by - amitb.UNKNOWN (DESKTOP-GIFQ7HQ)
//          at - 13:33:56 15/12/2018
//
// using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
//

`resetall
`timescale 1ns/10ps
module Checker#(
  parameter Amba_Word = 24,
  parameter Amba_Addr_Depth = 13,
  parameter Weight_precision = 5
)
(
  cat_recognizer_interface.checkr_coveragr checker_Interface
);

integer  clocks_counter=0;

  property reset_active;
            @( checker_Interface.rst) (checker_Interface.rst==1) |-> (checker_Interface.CatRecOut!=1);
  endproperty

  assert property(reset_active)
  else $error("problem with reset");
  cover property (reset_active);
  
  always @(posedge checker_Interface.clk)
  begin
  clocks_counter = clocks_counter + 1;
  end
  
  
	
	
endmodule
